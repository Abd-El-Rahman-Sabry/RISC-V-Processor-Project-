// RISC-V Core Implementation
// Authors: Abd-El-Rahman Sabry, Mahmoud Ahmed Mahmoud Abd-El-Halim
// Date: September 2024
// Description: This module implements a basic RISC-V processor core, including
// the instruction fetch, decode, execute, memory access, and write-back stages.
//
// Copyright (c) 2024 Abd-El-Rahman Sabry, Mahmoud Ahmed Mahmoud Abd-El-Halim
// All rights reserved.
// 
// This source code is proprietary and may not be reproduced, distributed,
// or transmitted in any form or by any means without the prior written
// permission of the authors.

`timescale 1ns/1ps



module tb;
    

    initial begin
        
        $display("Welcome to the RISC V Project."); 
        $display("Welcome to the RISC V Project."); 
        
        $finish; 
    end

endmodule